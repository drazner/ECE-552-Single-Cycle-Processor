
module p4(clk, rst, ,write_en, rf1, rf1_out, rf2, rf2_out, pc, pc_out, dm, dm_out, alu, alu_out, instr, instr_out, D_compute, D_compute_out, D_compute_imm, D_compute_imm_out, D_lw, D_lw_out, D_sw, D_sw_out, D_lhb, D_lhb_out,
		D_llb, D_llb_out, D_b, D_b_out, D_br, D_br_out, D_pcs, D_pcs_out, D_hlt, D_hlt_out);

input clk, rst, write_en;
input [15:0] instr, dm, alu, pc, rf1, rf2;
input D_compute, D_compute_imm, D_lw, D_sw, D_lhb, D_llb, D_b, D_br, D_pcs, D_hlt;
output [15:0] instr_out, dm_out, alu_out, pc_out, rf1_out, rf2_out;
output D_compute_out, D_compute_imm_out, D_lw_out, D_sw_out, D_lhb_out, D_llb_out, D_b_out, D_br_out, D_pcs_out, D_hlt_out;

//rf1
dff rf1_0(.q(rf1_out[0]), .d(rf1[0]), .wen(write_en), .clk(clk), .rst(rst));
dff rf1_1(.q(rf1_out[1]), .d(rf1[1]), .wen(write_en), .clk(clk), .rst(rst));
dff rf1_2(.q(rf1_out[2]), .d(rf1[2]), .wen(write_en), .clk(clk), .rst(rst));
dff rf1_3(.q(rf1_out[3]), .d(rf1[3]), .wen(write_en), .clk(clk), .rst(rst));
dff rf1_4(.q(rf1_out[4]), .d(rf1[4]), .wen(write_en), .clk(clk), .rst(rst));
dff rf1_5(.q(rf1_out[5]), .d(rf1[5]), .wen(write_en), .clk(clk), .rst(rst));
dff rf1_6(.q(rf1_out[6]), .d(rf1[6]), .wen(write_en), .clk(clk), .rst(rst));
dff rf1_7(.q(rf1_out[7]), .d(rf1[7]), .wen(write_en), .clk(clk), .rst(rst));
dff rf1_8(.q(rf1_out[8]), .d(rf1[8]), .wen(write_en), .clk(clk), .rst(rst));
dff rf1_9(.q(rf1_out[9]), .d(rf1[9]), .wen(write_en), .clk(clk), .rst(rst));
dff rf1_10(.q(rf1_out[10]), .d(rf1[10]), .wen(write_en), .clk(clk), .rst(rst));
dff rf1_11(.q(rf1_out[11]), .d(rf1[11]), .wen(write_en), .clk(clk), .rst(rst));
dff rf1_12(.q(rf1_out[12]), .d(rf1[12]), .wen(write_en), .clk(clk), .rst(rst));
dff rf1_13(.q(rf1_out[13]), .d(rf1[13]), .wen(write_en), .clk(clk), .rst(rst));
dff rf1_14(.q(rf1_out[14]), .d(rf1[14]), .wen(write_en), .clk(clk), .rst(rst));
dff rf1_15(.q(rf1_out[15]), .d(rf1[15]), .wen(write_en), .clk(clk), .rst(rst));

//rf2
dff rf2_0(.q(rf2_out[0]), .d(rf2[0]), .wen(write_en), .clk(clk), .rst(rst));
dff rf2_1(.q(rf2_out[1]), .d(rf2[1]), .wen(write_en), .clk(clk), .rst(rst));
dff rf2_2(.q(rf2_out[2]), .d(rf2[2]), .wen(write_en), .clk(clk), .rst(rst));
dff rf2_3(.q(rf2_out[3]), .d(rf2[3]), .wen(write_en), .clk(clk), .rst(rst));
dff rf2_4(.q(rf2_out[4]), .d(rf2[4]), .wen(write_en), .clk(clk), .rst(rst));
dff rf2_5(.q(rf2_out[5]), .d(rf2[5]), .wen(write_en), .clk(clk), .rst(rst));
dff rf2_6(.q(rf2_out[6]), .d(rf2[6]), .wen(write_en), .clk(clk), .rst(rst));
dff rf2_7(.q(rf2_out[7]), .d(rf2[7]), .wen(write_en), .clk(clk), .rst(rst));
dff rf2_8(.q(rf2_out[8]), .d(rf2[8]), .wen(write_en), .clk(clk), .rst(rst));
dff rf2_9(.q(rf2_out[9]), .d(rf2[9]), .wen(write_en), .clk(clk), .rst(rst));
dff rf2_10(.q(rf2_out[10]), .d(rf2[10]), .wen(write_en), .clk(clk), .rst(rst));
dff rf2_11(.q(rf2_out[11]), .d(rf2[11]), .wen(write_en), .clk(clk), .rst(rst));
dff rf2_12(.q(rf2_out[12]), .d(rf2[12]), .wen(write_en), .clk(clk), .rst(rst));
dff rf2_13(.q(rf2_out[13]), .d(rf2[13]), .wen(write_en), .clk(clk), .rst(rst));
dff rf2_14(.q(rf2_out[14]), .d(rf2[14]), .wen(write_en), .clk(clk), .rst(rst));
dff rf2_15(.q(rf2_out[15]), .d(rf2[15]), .wen(write_en), .clk(clk), .rst(rst));

//pc
dff pc_dff0(.q(pc_out[0]), .d(pc[0]), .wen(write_en), .clk(clk), .rst(rst));
dff pc_dff1(.q(pc_out[1]), .d(pc[1]), .wen(write_en), .clk(clk), .rst(rst));
dff pc_dff2(.q(pc_out[2]), .d(pc[2]), .wen(write_en), .clk(clk), .rst(rst));
dff pc_dff3(.q(pc_out[3]), .d(pc[3]), .wen(write_en), .clk(clk), .rst(rst));
dff pc_dff4(.q(pc_out[4]), .d(pc[4]), .wen(write_en), .clk(clk), .rst(rst));
dff pc_dff5(.q(pc_out[5]), .d(pc[5]), .wen(write_en), .clk(clk), .rst(rst));
dff pc_dff6(.q(pc_out[6]), .d(pc[6]), .wen(write_en), .clk(clk), .rst(rst));
dff pc_dff7(.q(pc_out[7]), .d(pc[7]), .wen(write_en), .clk(clk), .rst(rst));
dff pc_dff8(.q(pc_out[8]), .d(pc[8]), .wen(write_en), .clk(clk), .rst(rst));
dff pc_dff9(.q(pc_out[9]), .d(pc[9]), .wen(write_en), .clk(clk), .rst(rst));
dff pc_dff10(.q(pc_out[10]), .d(pc[10]), .wen(write_en), .clk(clk), .rst(rst));
dff pc_dff11(.q(pc_out[11]), .d(pc[11]), .wen(write_en), .clk(clk), .rst(rst));
dff pc_dff12(.q(pc_out[12]), .d(pc[12]), .wen(write_en), .clk(clk), .rst(rst));
dff pc_dff13(.q(pc_out[13]), .d(pc[13]), .wen(write_en), .clk(clk), .rst(rst));
dff pc_dff14(.q(pc_out[14]), .d(pc[14]), .wen(write_en), .clk(clk), .rst(rst));
dff pc_dff15(.q(pc_out[15]), .d(pc[15]), .wen(write_en), .clk(clk), .rst(rst));

//alu
dff alu0(.q(alu_out[0]), .d(alu[0]), .wen(write_en), .clk(clk), .rst(rst));
dff alu1(.q(alu_out[1]), .d(alu[1]), .wen(write_en), .clk(clk), .rst(rst));
dff alu2(.q(alu_out[2]), .d(alu[2]), .wen(write_en), .clk(clk), .rst(rst));
dff alu3(.q(alu_out[3]), .d(alu[3]), .wen(write_en), .clk(clk), .rst(rst));
dff alu4(.q(alu_out[4]), .d(alu[4]), .wen(write_en), .clk(clk), .rst(rst));
dff alu5(.q(alu_out[5]), .d(alu[5]), .wen(write_en), .clk(clk), .rst(rst));
dff alu6(.q(alu_out[6]), .d(alu[6]), .wen(write_en), .clk(clk), .rst(rst));
dff alu7(.q(alu_out[7]), .d(alu[7]), .wen(write_en), .clk(clk), .rst(rst));
dff alu8(.q(alu_out[8]), .d(alu[8]), .wen(write_en), .clk(clk), .rst(rst));
dff alu9(.q(alu_out[9]), .d(alu[9]), .wen(write_en), .clk(clk), .rst(rst));
dff alu10(.q(alu_out[10]), .d(alu[10]), .wen(write_en), .clk(clk), .rst(rst));
dff alu11(.q(alu_out[11]), .d(alu[11]), .wen(write_en), .clk(clk), .rst(rst));
dff alu12(.q(alu_out[12]), .d(alu[12]), .wen(write_en), .clk(clk), .rst(rst));
dff alu13(.q(alu_out[13]), .d(alu[13]), .wen(write_en), .clk(clk), .rst(rst));
dff alu14(.q(alu_out[14]), .d(alu[14]), .wen(write_en), .clk(clk), .rst(rst));
dff alu15(.q(alu_out[15]), .d(alu[15]), .wen(write_en), .clk(clk), .rst(rst));


//dm
dff dm0(.q(dm_out[0]), .d(dm[0]), .wen(write_en), .clk(clk), .rst(rst));
dff dm1(.q(dm_out[1]), .d(dm[1]), .wen(write_en), .clk(clk), .rst(rst));
dff dm2(.q(dm_out[2]), .d(dm[2]), .wen(write_en), .clk(clk), .rst(rst));
dff dm3(.q(dm_out[3]), .d(dm[3]), .wen(write_en), .clk(clk), .rst(rst));
dff dm4(.q(dm_out[4]), .d(dm[4]), .wen(write_en), .clk(clk), .rst(rst));
dff dm5(.q(dm_out[5]), .d(dm[5]), .wen(write_en), .clk(clk), .rst(rst));
dff dm6(.q(dm_out[6]), .d(dm[6]), .wen(write_en), .clk(clk), .rst(rst));
dff dm7(.q(dm_out[7]), .d(dm[7]), .wen(write_en), .clk(clk), .rst(rst));
dff dm8(.q(dm_out[8]), .d(dm[8]), .wen(write_en), .clk(clk), .rst(rst));
dff dm9(.q(dm_out[9]), .d(dm[9]), .wen(write_en), .clk(clk), .rst(rst));
dff dm10(.q(dm_out[10]), .d(dm[10]), .wen(write_en), .clk(clk), .rst(rst));
dff dm11(.q(dm_out[11]), .d(dm[11]), .wen(write_en), .clk(clk), .rst(rst));
dff dm12(.q(dm_out[12]), .d(dm[12]), .wen(write_en), .clk(clk), .rst(rst));
dff dm13(.q(dm_out[13]), .d(dm[13]), .wen(write_en), .clk(clk), .rst(rst));
dff dm14(.q(dm_out[14]), .d(dm[14]), .wen(write_en), .clk(clk), .rst(rst));
dff dm15(.q(dm_out[15]), .d(dm[15]), .wen(write_en), .clk(clk), .rst(rst));

//instr
dff instr_dff0(.q(instr_out[0]), .d(instr[0]), .wen(write_en), .clk(clk), .rst(rst));
dff instr_dff1(.q(instr_out[1]), .d(instr[1]), .wen(write_en), .clk(clk), .rst(rst));
dff instr_dff2(.q(instr_out[2]), .d(instr[2]), .wen(write_en), .clk(clk), .rst(rst));
dff instr_dff3(.q(instr_out[3]), .d(instr[3]), .wen(write_en), .clk(clk), .rst(rst));
dff instr_dff4(.q(instr_out[4]), .d(instr[4]), .wen(write_en), .clk(clk), .rst(rst));
dff instr_dff5(.q(instr_out[5]), .d(instr[5]), .wen(write_en), .clk(clk), .rst(rst));
dff instr_dff6(.q(instr_out[6]), .d(instr[6]), .wen(write_en), .clk(clk), .rst(rst));
dff instr_dff7(.q(instr_out[7]), .d(instr[7]), .wen(write_en), .clk(clk), .rst(rst));
dff instr_dff8(.q(instr_out[8]), .d(instr[8]), .wen(write_en), .clk(clk), .rst(rst));
dff instr_dff9(.q(instr_out[9]), .d(instr[9]), .wen(write_en), .clk(clk), .rst(rst));
dff instr_dff10(.q(instr_out[10]), .d(instr[10]), .wen(write_en), .clk(clk), .rst(rst));
dff instr_dff11(.q(instr_out[11]), .d(instr[11]), .wen(write_en), .clk(clk), .rst(rst));
dff instr_dff12(.q(instr_out[12]), .d(instr[12]), .wen(write_en), .clk(clk), .rst(rst));
dff instr_dff13(.q(instr_out[13]), .d(instr[13]), .wen(write_en), .clk(clk), .rst(rst));
dff instr_dff14(.q(instr_out[14]), .d(instr[14]), .wen(write_en), .clk(clk), .rst(rst));
dff instr_dff15(.q(instr_out[15]), .d(instr[15]), .wen(write_en), .clk(clk), .rst(rst));



//DECODE SIGNALS
dff D_compute_dff(.q(D_compute_out), .d(D_compute), .wen(write_en), .clk(clk), .rst(rst));
dff D_compute_imm_dff(.q(D_compute_imm_out), .d(D_compute_imm), .wen(write_en), .clk(clk), .rst(rst));
dff D_lw_dff(.q(D_lw_out), .d(D_lw), .wen(write_en), .clk(clk), .rst(rst));
dff D_sw_dff(.q(D_sw_out), .d(D_sw), .wen(write_en), .clk(clk), .rst(rst));
dff D_lhb_dff(.q(D_lhb_out), .d(D_lhb), .wen(write_en), .clk(clk), .rst(rst));
dff D_llb_dff(.q(D_llb_out), .d(D_llb), .wen(write_en), .clk(clk), .rst(rst));
dff D_b_dff(.q(D_b_out), .d(D_b), .wen(write_en), .clk(clk), .rst(rst));
dff D_br_dff(.q(D_br_out), .d(D_br), .wen(write_en), .clk(clk), .rst(rst));
dff D_pcs_dff(.q(D_pcs_out), .d(D_pcs), .wen(write_en), .clk(clk), .rst(rst));
dff D_hlt_dff(.q(D_hlt_out), .d(D_hlt), .wen(write_en), .clk(clk), .rst(rst));






endmodule