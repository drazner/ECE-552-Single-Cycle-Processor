
module ROR(result, A, imm); 

//16 bit input reg,4 bit immediate
input[15:0] A;
input[3:0] imm;

//16 bit output
output[15:0] result;

assign result = (imm == 4'b0000) ? A[15:0]:
		(imm == 4'b0001) ? {A[0],A[15:1]}:
		(imm == 4'b0010) ? {A[1:0],A[15:2]}:
		(imm == 4'b0011) ? {A[2:0],A[15:3]}:
		(imm == 4'b0100) ? {A[3:0],A[15:4]}:
		(imm == 4'b0101) ? {A[4:0],A[15:5]}:
		(imm == 4'b0110) ? {A[5:0],A[15:6]}:
		(imm == 4'b0111) ? {A[6:0],A[15:7]}:
		(imm == 4'b1000) ? {A[7:0],A[15:8]}:
		(imm == 4'b1001) ? {A[8:0],A[15:9]}:
		(imm == 4'b1010) ? {A[9:0],A[15:10]}:
		(imm == 4'b1010) ? {A[10:0],A[15:11]}:
		(imm == 4'b1100) ? {A[11:0],A[15:12]}:
		(imm == 4'b1101) ? {A[12:0],A[15:13]}:
		(imm == 4'b1110) ? {A[13:0],A[15:14]}:
		(imm == 4'b1111) ? {A[14:0],A[15]}:
		A[15:0]; 
		




endmodule
